module not_32bit(output [31:0] result, input [31:0] a);

	not_1bit not0 (result[0], a[0]);
	not_1bit not1 (result[1], a[1]);
	not_1bit not2 (result[2], a[2]);
	not_1bit not3 (result[3], a[3]);
	not_1bit not4 (result[4], a[4]);
	not_1bit not5 (result[5], a[5]);
	not_1bit not6 (result[6], a[6]);
	not_1bit not7 (result[7], a[7]);
	not_1bit not8 (result[8], a[8]);
	not_1bit not9 (result[9], a[9]);
	not_1bit not10 (result[10], a[10]);
	not_1bit not11 (result[11], a[11]);
	not_1bit not12 (result[12], a[12]);
	not_1bit not13 (result[13], a[13]);
	not_1bit not14 (result[14], a[14]);
	not_1bit not15 (result[15], a[15]);
	not_1bit not16 (result[16], a[16]);
	not_1bit not17 (result[17], a[17]);
	not_1bit not18 (result[18], a[18]);
	not_1bit not19 (result[19], a[19]);
	not_1bit not20 (result[20], a[20]);
	not_1bit not21 (result[21], a[21]);
	not_1bit not22 (result[22], a[22]);
	not_1bit not23 (result[23], a[23]);
	not_1bit not24 (result[24], a[24]);
	not_1bit not25 (result[25], a[25]);
	not_1bit not26 (result[26], a[26]);
	not_1bit not27 (result[27], a[27]);
	not_1bit not28 (result[28], a[28]);
	not_1bit not29 (result[29], a[29]);
	not_1bit not30 (result[30], a[30]);
	not_1bit not31 (result[31], a[31]);


endmodule