module not_1bit(output result, input a);

	not not1(result, a);

endmodule